Amplitude Response of Chebyshev Filter

V1 in 0 dc 0 ac 1
R0 in 1 1
C1 1 0 4.43m ic=0
L2 1 2 3.16m
C3 2 0 6.28m ic=0
L4 2 3 2.23m
RL 3 0 1.9841

.control
ac dec 10 1 1000
wrdata resp_cheby.txt vdb(3)
.endc

.end